package pseudo_rand_num_gen_pkg;
typedef enum logic[1:0] {
    RESET   = 2'b00,
    RUN     = 2'b01,
    DONE    = 2'b10,
    STATEX  = 2'bxx
} st_prng_state;
endpackage
